//localparam MAX_CLKS = 1000000;

localparam BLANK     = 3'd0;
localparam LIME      = 3'd1;
localparam ORANGE    = 3'd2;
localparam GRAPE     = 3'd3;
localparam BANANA    = 3'd4;
localparam BLUEBERRY = 3'd5;
localparam CHERRY    = 3'd6;
localparam COCONUT   = 3'd7;

